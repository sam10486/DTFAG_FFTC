`ifndef DEFINE_SVH
`define DEFINE_SVH

`timescale 10ns / 1ps
`define D_width 64
`define doulbe_D_width 128
`define radix_r 16
`define radix_width 4 //log2(radix)
`define ROMA_width 6


`endif 